library ieee;
use ieee.std_logic_1164.all;

entity ClkDivider is 
	port(clk : in std_logic;
			)